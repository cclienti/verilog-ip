//                              -*- Mode: Verilog -*-
// Filename        : cmpgt_tb.v
// Description     : Signed-unsigned dual-mode comparator testbench
// Author          : Christophe Clienti
// Created On      : Wed Feb 16 15:47:14 2013
// Last Modified By: Christophe Clienti
// Last Modified On: Wed Feb 16 15:47:14 2013
// Update Count    : 0
// Status          : Unknown, Use with caution!
// Copyright (C) 2013-2016 Christophe Clienti - All Rights Reserved

`timescale 1 ns / 100 ps

module cmpgt_tb () ;
   parameter WIDTH = 16;

   reg [WIDTH-1:0] a, b;
   reg             is_signed;
   wire            out;

   integer         cpt;


   cmpgt #(.WIDTH(WIDTH))
   DUT(.out(out), .is_signed(is_signed), .a(a), .b(b));


   initial  begin
      $dumpfile ("cmpgt_tb.vcd");
      $dumpvars;
   end


   initial begin
      cpt = 0;
      #1000 $finish;
   end


   always
     #2 cpt <= cpt + 1;


   always @ (cpt)
     begin
        case (cpt)
          0: begin
             a <= 0;
             b <= 0;
             is_signed <= 0;
          end
          1: begin
             a <= -1;
             b <= 1;
             is_signed <= 0;
          end
          2: begin
             a <= -1;
             b <= 1;
             is_signed <= 1;
          end
          3: begin
             a = 2;
             b = -1;
             is_signed = 0;
          end
          4: begin
             a = 2;
             b = -1;
             is_signed = 1;
          end
          5: begin
             a = 2;
             b = 1;
             is_signed = 0;
          end
          6: begin
             a = 2;
             b = 1;
             is_signed = 1;
          end
          7: begin
             a = 1;
             b = 2;
             is_signed = 0;
          end
          8: begin
             a = 1;
             b = 2;
             is_signed = 1;
          end
          9: begin
             a = -2;
             b = -1;
             is_signed = 1;
          end
          10: begin
             a = -2;
             b = -1;
             is_signed = 0;
          end
          11: begin
             a = -1;
             b = -2;
             is_signed = 1;
          end
          12: begin
             a = -1;
             b = -2;
             is_signed = 0;
          end
          13: $finish;

        endcase // case (cpt)
     end

endmodule // cmpgt_tb
